library ieee;
use ieee.std_logic_1164.all;

entity top_level is
    port(

        

    );
end top_level;