--in every project there will always be a library declared by default, implicitly: the work library
--it can be used by every file of your project in any level so that every structure you make can be used anywhere

--any library is gonna contain a number of packages

library ieee;
use ieee.std_logic_1164.all; --the "all" means we are gonna use all of the package (std_logic_1164)