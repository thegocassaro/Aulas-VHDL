library ieee;
use ieee.std_logic_1164.all;

entity prio_encoder32 is

    port(
        r: in std_logic_vector(2 downto 0);
        code: out std_logic_vector(1 downto 0)
        );

end prio_encoder32;


architecture cond_arch of prio_encoder32 is

begin
    code <= "11" when (r(2)='1') else
            "10" when (r(1)='1') else
            "01" when (r(0)='1') else
            "00";

end cond_arch;