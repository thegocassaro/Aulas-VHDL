entity TESTE_01 is 
end entity;

architecture sim of TESTE_01 is

begin

    process is
    begin

        report "Hello World!";
        wait;

    end process;

end architecture;